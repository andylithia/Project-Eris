module CTC (
	//input			cph1,
	input			cph2,
	input			pon,
	input			is,
	input			carry
	output			ws,
	output			sync,

	output [7:0]	kr,
	input [4:0]		kc
);




endmodule // CTC